----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:17:31 05/04/2022 
-- Design Name: 
-- Module Name:    ROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- 16x8 ROM
-- IVH -> lectures -> 07 -> slide 76
entity ROM is
port (
		ADDRESS : in integer range 0 to 1000;
		DATA : out std_logic_vector(127 downto 0);
		CLK : in std_logic
		);
end ROM;

architecture rtl of ROM is
	type rom_array is array (0 to 57) of std_logic_vector(127 downto 0);
	constant rom: rom_array := (
										-- LEFT 1
										"01111111010001010100010101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --11	--1
										"00000000011111110100010101000101011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --10	--2
										"00000000000000000111111101000101010001010111111100000000000000000000000000000000000000000000000000000000000000000000000000000000", --7	--3
										
										"00000000000000000000000001111111010001010100010101111111000000000000000000000000000000000000000000000000000000000000000000000000", --6	--4
										"00000000000000000000000000000000011111110100010101000101011111110000000000000000000000000000000000000000000000000000000000000000", --3	--5
										"00000000000000000000000000000000000000000111111101000101010001010111111100000000000000000000000000000000000000000000000000000000", --2	--6
										
										"00000000000000000000000000000000000000000000000001111111010001010100010101111111000000000000000000000000000000000000000000000000", --13	--7
										"00000000000000000000000000000000000000000000000000000000011111110100010101000101011111110000000000000000000000000000000000000000", --12	--8
										"00000000000000000000000000000000000000000000000000000000000000000111111101000101010001010111111100000000000000000000000000000000", --9	--9
										
										"00000000000000000000000000000000000000000000000000000000000000000000000001111111010001010100010101111111000000000000000000000000", --8	--10
										"00000000000000000000000000000000000000000000000000000000000000000000000000000000011111110100010101000101011111110000000000000000", --5	--11
										"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101000101010001010111111100000000", --4	--12
										"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111010001010100010101111111", --1	--13
										
										-- RIGHT 1
										"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111010001010100010101111111", --1	--13
										"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101000101010001010111111100000000", --4	--12
										"00000000000000000000000000000000000000000000000000000000000000000000000000000000011111110100010101000101011111110000000000000000", --5	--11
										"00000000000000000000000000000000000000000000000000000000000000000000000001111111010001010100010101111111000000000000000000000000", --8	--10
										
										"00000000000000000000000000000000000000000000000000000000000000000111111101000101010001010111111100000000000000000000000000000000", --9	--9
										"00000000000000000000000000000000000000000000000000000000011111110100010101000101011111110000000000000000000000000000000000000000", --12	--8
										"00000000000000000000000000000000000000000000000001111111010001010100010101111111000000000000000000000000000000000000000000000000", --13	--7
										"00000000000000000000000000000000000000000111111101000101010001010111111100000000000000000000000000000000000000000000000000000000", --2	--6
										"00000000000000000000000000000000011111110100010101000101011111110000000000000000000000000000000000000000000000000000000000000000", --3	--5
										"00000000000000000000000001111111010001010100010101111111000000000000000000000000000000000000000000000000000000000000000000000000", --6	--4
										"00000000000000000111111101000101010001010111111100000000000000000000000000000000000000000000000000000000000000000000000000000000", --7	--3
										"00000000011111110100010101000101011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --10	--2
										"01111111010001010100010101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --11	--1
										
										-- LEFT 2
										"01111111010001010100010101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --11	--1
										"00000000011111110100010101000101011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --10	--2
										"00000000000000000111111101000101010001010111111100000000000000000000000000000000000000000000000000000000000000000000000000000000", --7	--3
										
										"00000000000000000000000001111111010001010100010101111111000000000000000000000000000000000000000000000000000000000000000000000000", --6	--4
										"00000000000000000000000000000000011111110100010101000101011111110000000000000000000000000000000000000000000000000000000000000000", --3	--5
										"00000000000000000000000000000000000000000111111101000101010001010111111100000000000000000000000000000000000000000000000000000000", --2	--6
										
										"00000000000000000000000000000000000000000000000001111111010001010100010101111111000000000000000000000000000000000000000000000000", --13	--7
										"00000000000000000000000000000000000000000000000000000000011111110100010101000101011111110000000000000000000000000000000000000000", --12	--8
										"00000000000000000000000000000000000000000000000000000000000000000111111101000101010001010111111100000000000000000000000000000000", --9	--9
										
										"00000000000000000000000000000000000000000000000000000000000000000000000001111111010001010100010101111111000000000000000000000000", --8	--10
										"00000000000000000000000000000000000000000000000000000000000000000000000000000000011111110100010101000101011111110000000000000000", --5	--11
										"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101000101010001010111111100000000", --4	--12
										"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111010001010100010101111111", --1	--13
										
										-- RIGHT 2
										"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111010001010100010101111111", --1	--13
										"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101000101010001010111111100000000", --4	--12
										"00000000000000000000000000000000000000000000000000000000000000000000000000000000011111110100010101000101011111110000000000000000", --5	--11
										"00000000000000000000000000000000000000000000000000000000000000000000000001111111010001010100010101111111000000000000000000000000", --8	--10
										
										"00000000000000000000000000000000000000000000000000000000000000000111111101000101010001010111111100000000000000000000000000000000", --9	--9
										"00000000000000000000000000000000000000000000000000000000011111110100010101000101011111110000000000000000000000000000000000000000", --12	--8
										"00000000000000000000000000000000000000000000000001111111010001010100010101111111000000000000000000000000000000000000000000000000", --13	--7
										"00000000000000000000000000000000000000000111111101000101010001010111111100000000000000000000000000000000000000000000000000000000", --2	--6
										"00000000000000000000000000000000011111110100010101000101011111110000000000000000000000000000000000000000000000000000000000000000", --3	--5
										"00000000000000000000000001111111010001010100010101111111000000000000000000000000000000000000000000000000000000000000000000000000", --6	--4
										"00000000000000000111111101000101010001010111111100000000000000000000000000000000000000000000000000000000000000000000000000000000", --7	--3
										"00000000011111110100010101000101011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --10	--2
										"01111111010001010100010101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --11	--1

										-- ANIMATION
										"01010101101010100101010110101010010101011010101001010101101010100101010110101010010101011010101001010101101010100101010110101010", --14
										"10101010010101011010101001010101101010100101010110101010010101011010101001010101101010100101010110101010010101011010101001010101", --15
										"01010101101010100101010110101010010101011010101001010101101010100101010110101010010101011010101001010101101010100101010110101010", --14
										"10101010010101011010101001010101101010100101010110101010010101011010101001010101101010100101010110101010010101011010101001010101", --15
										"01010101101010100101010110101010010101011010101001010101101010100101010110101010010101011010101001010101101010100101010110101010", --14
										"10101010010101011010101001010101101010100101010110101010010101011010101001010101101010100101010110101010010101011010101001010101" --15 -- 83
										);
begin
	result: process (ADDRESS) is
	begin
		--if (rising_edge(CLK) then
			DATA <= rom(ADDRESS);
		--end if;
	end process;
end architecture;

